module tabla01_SOP();

// Pruebas

// Ya hay algo que no quiero perder (quiero dejarlo guardado como una "versión" de mi código.



endmodule
