module tabla01_POS();





endmodule
