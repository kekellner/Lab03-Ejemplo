module tabla01_POS();

// Empezar todo mi código...

// pruebas

// más pruebas

// ya avancé algo significativo



endmodule
